module DFF
(
input clk,rst,
input signed[31:0] d,
output reg signed [31:0] q 
);
    
always@ (posedge clk, posedge rst)
    if(rst)
        q<=0;
    else
        q<=d;
endmodule
