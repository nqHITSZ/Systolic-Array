//process element
module mult
(
input 
)
